module vedic_16bit_mul (
    input [15:0] a,
    input [15:0] b,
    output [31:0] m
);

    wire [15:0] p0, p1, p2, p3; 
    
    wire [15:0] temp1, temp2, temp3; 
    wire cout1, cout2, cout3;
    wire cin3;

    vedic_8bit_mul m1 (.a(a[7:0]), .b(b[7:0]), .m(p0));
    vedic_8bit_mul m2 (.a(a[7:0]), .b(b[15:8]), .m(p1));
    vedic_8bit_mul m3 (.a(a[15:8]), .b(b[7:0]), .m(p2));
    vedic_8bit_mul m4 (.a(a[15:8]), .b(b[15:8]), .m(p3));

    cla_nbit #(.WIDTH(16)) adder1 (  
        .a(p1),
        .b(p2),
        .cin(1'b0),
        .sum(temp1),
        .cout(cout1)
    );

    cla_nbit #(.WIDTH(16)) adder2 (
        .a(temp1),
        .b({8'h00, p0[15:8]}),
        .cin(1'b0),
        .sum(temp2),
        .cout(cout2)
    );

    assign cin3 = cout1 | cout2;

    cla_nbit #(.WIDTH(16)) adder3 (
        .a({7'b0000000, cin3, temp2[15:8]}),  
        .b(p3),
        .cin(1'b0),
        .sum(temp3),
        .cout(cout3)
    );

    assign m = {temp3, temp2[7:0], p0[7:0]};

endmodule

/*
710     65407   65400   4277617800 (4277617800)
720     65407   65401   4277683207 (4277683207)
730     65407   65402   4277748614 (4277748614)
740     65407   65403   4277814021 (4277814021)
750     65407   65404   4277879428 (4277879428)
760     65407   65405   4277944835 (4277944835)
770     65407   65406   4278010242 (4278010242)
780     65407   65407   4278075649 (4278075649)
790     65407   65408   4278141056 (4278141056)
800     65407   65409   4278206463 (4278206463)
810     65408   65400   4277683200 (4277683200)
820     65408   65401   4277748608 (4277748608)
830     65408   65402   4277814016 (4277814016)
840     65408   65403   4277879424 (4277879424)
850     65408   65404   4277944832 (4277944832)
860     65408   65405   4278010240 (4278010240)
870     65408   65406   4278075648 (4278075648)
880     65408   65407   4278141056 (4278141056)
890     65408   65408   4278206464 (4278206464)
900     65408   65409   4278271872 (4278271872)
910     65409   65400   4277748600 (4277748600)
920     65409   65401   4277814009 (4277814009)
930     65409   65402   4277879418 (4277879418)
940     65409   65403   4277944827 (4277944827)
950     65409   65404   4278010236 (4278010236)
960     65409   65405   4278075645 (4278075645)
970     65409   65406   4278141054 (4278141054)
980     65409   65407   4278206463 (4278206463)
990     65409   65408   4278271872 (4278271872)
1000    65409   65409   4278337281 (4278337281)
*/
